class stimulus;
  rand   logic[31:0]  valueA  ;
  rand   logic[31:0]  valueB  ;
  shortreal floatA = valueA;
  shortreal floatB = valueB;
  
  //constraint distribution {value dist { 0  := 1 , 1 := 1 }; } 
endclass
